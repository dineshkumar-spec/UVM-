interface intf;
  logic a,b;
  logic sum,carry;
endinterface
