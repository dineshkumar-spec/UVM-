interface intf;
  logic clk;
  logic reset;
  logic d;
  logic q;
endinterface
